`timescale 1ns/10ps

module ALU(input[3:0] OPCODE, input[7:0] R1, input[7:0] R2, output[7:0] ROUT);
endmodule
